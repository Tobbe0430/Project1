module IF_ID 	
(
	clk_i,
	inst_addr_i,
	inst_i,
	hd_i,
	flush_i,
	mux2_o,
	hd_o,
	op_o,
	inst_addr1_o,
	inst_addr2_o,
	rs1_o,
	rt1_o,
	rs2_o,
	rt2_o,
	sign16_o,
	rd_o
);

input			clk_i;
input	[31:0]	inst_addr_i,inst_i;
input			hd_i,flush_i;
output	[25:0]	mux2_o;
output	??		hd_o;
output	[5:0]	op_o;
output	[31:0]	inst_addr1_o,inst_addr2_o;
output	[4:0]	rs1_o,rt1_o, rs2_o, rt2_o, rd_o;
output	[15:0]	sign16_o;

assign mux2_o = inst_i[25:0];
assign hd_o = ??
assign op_o = inst_i[5:0];
assign inst_addr1_o = inst_addr_i;
assign inst_addr2_o = inst_addr_i;
assign rs1_o = inst_i[25:21];
assign rs2_o = inst_i[25:21];
assign rt1_o = inst_i[20:16];
assign rt2_o = inst_i[20:16];
assign sign16_o = inst_i[15:0];
assign rd_o = inst_i[15:11];

reg 	[31:0] 	inst_addr;
reg 	[31:0]  inst;

WHAT ABOUT FLUSH THOUGH??????

always@(posedge clk_i) begin
    if(NO FLUSH MAYBE?)
        inst_addr <= inst_addr_i;
		inst <= inst_i;
end

endmodule 