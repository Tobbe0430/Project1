module Flush
(
	jump_i;
	branch_i;
	flush_o;
);

input	jump_i,branch_i;
output	flush_o;

endmodule